
module router4x144 (
    

    i_data0, i_data1, i_data2, i_data3, 
   

    o_val
 
);

  

  input[23:0] i_data0, i_data1, i_data2, i_data3;
  


  output [20*144 - 1 : 0 ] o_val;

  
  wire [143:0] select0, select1, select2, select3; 

  

  sel1x144 u_sel1x144_0 (.x_cor(i_data0[23:20]), .y_cor(i_data0[19:16]), .select(select0));
  sel1x144 u_sel1x144_1 (.x_cor(i_data1[23:20]), .y_cor(i_data1[19:16]), .select(select1));
  sel1x144 u_sel1x144_2 (.x_cor(i_data2[23:20]), .y_cor(i_data2[19:16]), .select(select2));
  sel1x144 u_sel1x144_3 (.x_cor(i_data3[23:20]), .y_cor(i_data3[19:16]), .select(select3));
  
addertree u_addertree_0 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[0], select2[0], select1[0], select0[0]}), .o_val(o_val[19:0]));
addertree u_addertree_1 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[1], select2[1], select1[1], select0[1]}), .o_val(o_val[39:20]));
addertree u_addertree_2 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[2], select2[2], select1[2], select0[2]}), .o_val(o_val[59:40]));
addertree u_addertree_3 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[3], select2[3], select1[3], select0[3]}), .o_val(o_val[79:60]));
addertree u_addertree_4 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[4], select2[4], select1[4], select0[4]}), .o_val(o_val[99:80]));
addertree u_addertree_5 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[5], select2[5], select1[5], select0[5]}), .o_val(o_val[119:100]));
addertree u_addertree_6 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[6], select2[6], select1[6], select0[6]}), .o_val(o_val[139:120]));
addertree u_addertree_7 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[7], select2[7], select1[7], select0[7]}), .o_val(o_val[159:140]));
addertree u_addertree_8 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[8], select2[8], select1[8], select0[8]}), .o_val(o_val[179:160]));
addertree u_addertree_9 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[9], select2[9], select1[9], select0[9]}), .o_val(o_val[199:180]));
addertree u_addertree_10 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[10], select2[10], select1[10], select0[10]}), .o_val(o_val[219:200]));
addertree u_addertree_11 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[11], select2[11], select1[11], select0[11]}), .o_val(o_val[239:220]));
addertree u_addertree_12 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[12], select2[12], select1[12], select0[12]}), .o_val(o_val[259:240]));
addertree u_addertree_13 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[13], select2[13], select1[13], select0[13]}), .o_val(o_val[279:260]));
addertree u_addertree_14 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[14], select2[14], select1[14], select0[14]}), .o_val(o_val[299:280]));
addertree u_addertree_15 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[15], select2[15], select1[15], select0[15]}), .o_val(o_val[319:300]));
addertree u_addertree_16 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[16], select2[16], select1[16], select0[16]}), .o_val(o_val[339:320]));
addertree u_addertree_17 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[17], select2[17], select1[17], select0[17]}), .o_val(o_val[359:340]));
addertree u_addertree_18 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[18], select2[18], select1[18], select0[18]}), .o_val(o_val[379:360]));
addertree u_addertree_19 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[19], select2[19], select1[19], select0[19]}), .o_val(o_val[399:380]));
addertree u_addertree_20 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[20], select2[20], select1[20], select0[20]}), .o_val(o_val[419:400]));
addertree u_addertree_21 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[21], select2[21], select1[21], select0[21]}), .o_val(o_val[439:420]));
addertree u_addertree_22 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[22], select2[22], select1[22], select0[22]}), .o_val(o_val[459:440]));
addertree u_addertree_23 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[23], select2[23], select1[23], select0[23]}), .o_val(o_val[479:460]));
addertree u_addertree_24 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[24], select2[24], select1[24], select0[24]}), .o_val(o_val[499:480]));
addertree u_addertree_25 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[25], select2[25], select1[25], select0[25]}), .o_val(o_val[519:500]));
addertree u_addertree_26 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[26], select2[26], select1[26], select0[26]}), .o_val(o_val[539:520]));
addertree u_addertree_27 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[27], select2[27], select1[27], select0[27]}), .o_val(o_val[559:540]));
addertree u_addertree_28 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[28], select2[28], select1[28], select0[28]}), .o_val(o_val[579:560]));
addertree u_addertree_29 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[29], select2[29], select1[29], select0[29]}), .o_val(o_val[599:580]));
addertree u_addertree_30 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[30], select2[30], select1[30], select0[30]}), .o_val(o_val[619:600]));
addertree u_addertree_31 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[31], select2[31], select1[31], select0[31]}), .o_val(o_val[639:620]));
addertree u_addertree_32 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[32], select2[32], select1[32], select0[32]}), .o_val(o_val[659:640]));
addertree u_addertree_33 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[33], select2[33], select1[33], select0[33]}), .o_val(o_val[679:660]));
addertree u_addertree_34 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[34], select2[34], select1[34], select0[34]}), .o_val(o_val[699:680]));
addertree u_addertree_35 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[35], select2[35], select1[35], select0[35]}), .o_val(o_val[719:700]));
addertree u_addertree_36 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[36], select2[36], select1[36], select0[36]}), .o_val(o_val[739:720]));
addertree u_addertree_37 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[37], select2[37], select1[37], select0[37]}), .o_val(o_val[759:740]));
addertree u_addertree_38 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[38], select2[38], select1[38], select0[38]}), .o_val(o_val[779:760]));
addertree u_addertree_39 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[39], select2[39], select1[39], select0[39]}), .o_val(o_val[799:780]));
addertree u_addertree_40 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[40], select2[40], select1[40], select0[40]}), .o_val(o_val[819:800]));
addertree u_addertree_41 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[41], select2[41], select1[41], select0[41]}), .o_val(o_val[839:820]));
addertree u_addertree_42 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[42], select2[42], select1[42], select0[42]}), .o_val(o_val[859:840]));
addertree u_addertree_43 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[43], select2[43], select1[43], select0[43]}), .o_val(o_val[879:860]));
addertree u_addertree_44 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[44], select2[44], select1[44], select0[44]}), .o_val(o_val[899:880]));
addertree u_addertree_45 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[45], select2[45], select1[45], select0[45]}), .o_val(o_val[919:900]));
addertree u_addertree_46 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[46], select2[46], select1[46], select0[46]}), .o_val(o_val[939:920]));
addertree u_addertree_47 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[47], select2[47], select1[47], select0[47]}), .o_val(o_val[959:940]));
addertree u_addertree_48 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[48], select2[48], select1[48], select0[48]}), .o_val(o_val[979:960]));
addertree u_addertree_49 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[49], select2[49], select1[49], select0[49]}), .o_val(o_val[999:980]));
addertree u_addertree_50 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[50], select2[50], select1[50], select0[50]}), .o_val(o_val[1019:1000]));
addertree u_addertree_51 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[51], select2[51], select1[51], select0[51]}), .o_val(o_val[1039:1020]));
addertree u_addertree_52 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[52], select2[52], select1[52], select0[52]}), .o_val(o_val[1059:1040]));
addertree u_addertree_53 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[53], select2[53], select1[53], select0[53]}), .o_val(o_val[1079:1060]));
addertree u_addertree_54 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[54], select2[54], select1[54], select0[54]}), .o_val(o_val[1099:1080]));
addertree u_addertree_55 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[55], select2[55], select1[55], select0[55]}), .o_val(o_val[1119:1100]));
addertree u_addertree_56 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[56], select2[56], select1[56], select0[56]}), .o_val(o_val[1139:1120]));
addertree u_addertree_57 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[57], select2[57], select1[57], select0[57]}), .o_val(o_val[1159:1140]));
addertree u_addertree_58 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[58], select2[58], select1[58], select0[58]}), .o_val(o_val[1179:1160]));
addertree u_addertree_59 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[59], select2[59], select1[59], select0[59]}), .o_val(o_val[1199:1180]));
addertree u_addertree_60 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[60], select2[60], select1[60], select0[60]}), .o_val(o_val[1219:1200]));
addertree u_addertree_61 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[61], select2[61], select1[61], select0[61]}), .o_val(o_val[1239:1220]));
addertree u_addertree_62 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[62], select2[62], select1[62], select0[62]}), .o_val(o_val[1259:1240]));
addertree u_addertree_63 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[63], select2[63], select1[63], select0[63]}), .o_val(o_val[1279:1260]));
addertree u_addertree_64 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[64], select2[64], select1[64], select0[64]}), .o_val(o_val[1299:1280]));
addertree u_addertree_65 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[65], select2[65], select1[65], select0[65]}), .o_val(o_val[1319:1300]));
addertree u_addertree_66 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[66], select2[66], select1[66], select0[66]}), .o_val(o_val[1339:1320]));
addertree u_addertree_67 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[67], select2[67], select1[67], select0[67]}), .o_val(o_val[1359:1340]));
addertree u_addertree_68 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[68], select2[68], select1[68], select0[68]}), .o_val(o_val[1379:1360]));
addertree u_addertree_69 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[69], select2[69], select1[69], select0[69]}), .o_val(o_val[1399:1380]));
addertree u_addertree_70 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[70], select2[70], select1[70], select0[70]}), .o_val(o_val[1419:1400]));
addertree u_addertree_71 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[71], select2[71], select1[71], select0[71]}), .o_val(o_val[1439:1420]));
addertree u_addertree_72 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[72], select2[72], select1[72], select0[72]}), .o_val(o_val[1459:1440]));
addertree u_addertree_73 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[73], select2[73], select1[73], select0[73]}), .o_val(o_val[1479:1460]));
addertree u_addertree_74 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[74], select2[74], select1[74], select0[74]}), .o_val(o_val[1499:1480]));
addertree u_addertree_75 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[75], select2[75], select1[75], select0[75]}), .o_val(o_val[1519:1500]));
addertree u_addertree_76 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[76], select2[76], select1[76], select0[76]}), .o_val(o_val[1539:1520]));
addertree u_addertree_77 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[77], select2[77], select1[77], select0[77]}), .o_val(o_val[1559:1540]));
addertree u_addertree_78 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[78], select2[78], select1[78], select0[78]}), .o_val(o_val[1579:1560]));
addertree u_addertree_79 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[79], select2[79], select1[79], select0[79]}), .o_val(o_val[1599:1580]));
addertree u_addertree_80 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[80], select2[80], select1[80], select0[80]}), .o_val(o_val[1619:1600]));
addertree u_addertree_81 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[81], select2[81], select1[81], select0[81]}), .o_val(o_val[1639:1620]));
addertree u_addertree_82 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[82], select2[82], select1[82], select0[82]}), .o_val(o_val[1659:1640]));
addertree u_addertree_83 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[83], select2[83], select1[83], select0[83]}), .o_val(o_val[1679:1660]));
addertree u_addertree_84 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[84], select2[84], select1[84], select0[84]}), .o_val(o_val[1699:1680]));
addertree u_addertree_85 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[85], select2[85], select1[85], select0[85]}), .o_val(o_val[1719:1700]));
addertree u_addertree_86 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[86], select2[86], select1[86], select0[86]}), .o_val(o_val[1739:1720]));
addertree u_addertree_87 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[87], select2[87], select1[87], select0[87]}), .o_val(o_val[1759:1740]));
addertree u_addertree_88 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[88], select2[88], select1[88], select0[88]}), .o_val(o_val[1779:1760]));
addertree u_addertree_89 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[89], select2[89], select1[89], select0[89]}), .o_val(o_val[1799:1780]));
addertree u_addertree_90 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[90], select2[90], select1[90], select0[90]}), .o_val(o_val[1819:1800]));
addertree u_addertree_91 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[91], select2[91], select1[91], select0[91]}), .o_val(o_val[1839:1820]));
addertree u_addertree_92 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[92], select2[92], select1[92], select0[92]}), .o_val(o_val[1859:1840]));
addertree u_addertree_93 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[93], select2[93], select1[93], select0[93]}), .o_val(o_val[1879:1860]));
addertree u_addertree_94 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[94], select2[94], select1[94], select0[94]}), .o_val(o_val[1899:1880]));
addertree u_addertree_95 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[95], select2[95], select1[95], select0[95]}), .o_val(o_val[1919:1900]));
addertree u_addertree_96 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[96], select2[96], select1[96], select0[96]}), .o_val(o_val[1939:1920]));
addertree u_addertree_97 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[97], select2[97], select1[97], select0[97]}), .o_val(o_val[1959:1940]));
addertree u_addertree_98 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[98], select2[98], select1[98], select0[98]}), .o_val(o_val[1979:1960]));
addertree u_addertree_99 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[99], select2[99], select1[99], select0[99]}), .o_val(o_val[1999:1980]));
addertree u_addertree_100 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[100], select2[100], select1[100], select0[100]}), .o_val(o_val[2019:2000]));
addertree u_addertree_101 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[101], select2[101], select1[101], select0[101]}), .o_val(o_val[2039:2020]));
addertree u_addertree_102 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[102], select2[102], select1[102], select0[102]}), .o_val(o_val[2059:2040]));
addertree u_addertree_103 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[103], select2[103], select1[103], select0[103]}), .o_val(o_val[2079:2060]));
addertree u_addertree_104 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[104], select2[104], select1[104], select0[104]}), .o_val(o_val[2099:2080]));
addertree u_addertree_105 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[105], select2[105], select1[105], select0[105]}), .o_val(o_val[2119:2100]));
addertree u_addertree_106 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[106], select2[106], select1[106], select0[106]}), .o_val(o_val[2139:2120]));
addertree u_addertree_107 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[107], select2[107], select1[107], select0[107]}), .o_val(o_val[2159:2140]));
addertree u_addertree_108 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[108], select2[108], select1[108], select0[108]}), .o_val(o_val[2179:2160]));
addertree u_addertree_109 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[109], select2[109], select1[109], select0[109]}), .o_val(o_val[2199:2180]));
addertree u_addertree_110 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[110], select2[110], select1[110], select0[110]}), .o_val(o_val[2219:2200]));
addertree u_addertree_111 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[111], select2[111], select1[111], select0[111]}), .o_val(o_val[2239:2220]));
addertree u_addertree_112 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[112], select2[112], select1[112], select0[112]}), .o_val(o_val[2259:2240]));
addertree u_addertree_113 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[113], select2[113], select1[113], select0[113]}), .o_val(o_val[2279:2260]));
addertree u_addertree_114 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[114], select2[114], select1[114], select0[114]}), .o_val(o_val[2299:2280]));
addertree u_addertree_115 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[115], select2[115], select1[115], select0[115]}), .o_val(o_val[2319:2300]));
addertree u_addertree_116 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[116], select2[116], select1[116], select0[116]}), .o_val(o_val[2339:2320]));
addertree u_addertree_117 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[117], select2[117], select1[117], select0[117]}), .o_val(o_val[2359:2340]));
addertree u_addertree_118 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[118], select2[118], select1[118], select0[118]}), .o_val(o_val[2379:2360]));
addertree u_addertree_119 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[119], select2[119], select1[119], select0[119]}), .o_val(o_val[2399:2380]));
addertree u_addertree_120 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[120], select2[120], select1[120], select0[120]}), .o_val(o_val[2419:2400]));
addertree u_addertree_121 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[121], select2[121], select1[121], select0[121]}), .o_val(o_val[2439:2420]));
addertree u_addertree_122 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[122], select2[122], select1[122], select0[122]}), .o_val(o_val[2459:2440]));
addertree u_addertree_123 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[123], select2[123], select1[123], select0[123]}), .o_val(o_val[2479:2460]));
addertree u_addertree_124 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[124], select2[124], select1[124], select0[124]}), .o_val(o_val[2499:2480]));
addertree u_addertree_125 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[125], select2[125], select1[125], select0[125]}), .o_val(o_val[2519:2500]));
addertree u_addertree_126 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[126], select2[126], select1[126], select0[126]}), .o_val(o_val[2539:2520]));
addertree u_addertree_127 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[127], select2[127], select1[127], select0[127]}), .o_val(o_val[2559:2540]));
addertree u_addertree_128 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[128], select2[128], select1[128], select0[128]}), .o_val(o_val[2579:2560]));
addertree u_addertree_129 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[129], select2[129], select1[129], select0[129]}), .o_val(o_val[2599:2580]));
addertree u_addertree_130 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[130], select2[130], select1[130], select0[130]}), .o_val(o_val[2619:2600]));
addertree u_addertree_131 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[131], select2[131], select1[131], select0[131]}), .o_val(o_val[2639:2620]));
addertree u_addertree_132 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[132], select2[132], select1[132], select0[132]}), .o_val(o_val[2659:2640]));
addertree u_addertree_133 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[133], select2[133], select1[133], select0[133]}), .o_val(o_val[2679:2660]));
addertree u_addertree_134 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[134], select2[134], select1[134], select0[134]}), .o_val(o_val[2699:2680]));
addertree u_addertree_135 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[135], select2[135], select1[135], select0[135]}), .o_val(o_val[2719:2700]));
addertree u_addertree_136 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[136], select2[136], select1[136], select0[136]}), .o_val(o_val[2739:2720]));
addertree u_addertree_137 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[137], select2[137], select1[137], select0[137]}), .o_val(o_val[2759:2740]));
addertree u_addertree_138 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[138], select2[138], select1[138], select0[138]}), .o_val(o_val[2779:2760]));
addertree u_addertree_139 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[139], select2[139], select1[139], select0[139]}), .o_val(o_val[2799:2780]));
addertree u_addertree_140 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[140], select2[140], select1[140], select0[140]}), .o_val(o_val[2819:2800]));
addertree u_addertree_141 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[141], select2[141], select1[141], select0[141]}), .o_val(o_val[2839:2820]));
addertree u_addertree_142 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[142], select2[142], select1[142], select0[142]}), .o_val(o_val[2859:2840]));
addertree u_addertree_143 (.i_val0(i_data0[15:0]), .i_val1(i_data1[15:0]), .i_val2(i_data2[15:0]), .i_val3(i_data3[15:0]), .sel({ select3[143], select2[143], select1[143], select0[143]}), .o_val(o_val[2879:2860]));

endmodule