module PPU(data_in, clk, en_encoder, en_pooling, row_size, index_pointer, row, data, out_port ,store, done);
    input[20 * 12 * 12 - 1 : 0] data_in;
    input clk, en_encoder, en_pooling;
    input [3:0] row_size;
    output[8 * 7 - 1 : 0] index_pointer;
    output[3 : 0] row;
    output[7 : 0] data;
    output store, done;
    output [31 : 0] out_port;
    
    wire [7 : 0] relu_out[0 : 143];
    wire [8 * 6 * 6 - 1 : 0] pooling_out;
    
    ReLU r0(.data_in(data_in[2879:2860]), .data_out(relu_out[0]));
    ReLU r1(.data_in(data_in[2859:2840]), .data_out(relu_out[1]));
    ReLU r2(.data_in(data_in[2839:2820]), .data_out(relu_out[2]));
    ReLU r3(.data_in(data_in[2819:2800]), .data_out(relu_out[3]));
    ReLU r4(.data_in(data_in[2799:2780]), .data_out(relu_out[4]));
    ReLU r5(.data_in(data_in[2779:2760]), .data_out(relu_out[5]));
    ReLU r6(.data_in(data_in[2759:2740]), .data_out(relu_out[6]));
    ReLU r7(.data_in(data_in[2739:2720]), .data_out(relu_out[7]));
    ReLU r8(.data_in(data_in[2719:2700]), .data_out(relu_out[8]));
    ReLU r9(.data_in(data_in[2699:2680]), .data_out(relu_out[9]));
    ReLU r10(.data_in(data_in[2679:2660]), .data_out(relu_out[10]));
    ReLU r11(.data_in(data_in[2659:2640]), .data_out(relu_out[11]));
    ReLU r12(.data_in(data_in[2639:2620]), .data_out(relu_out[12]));
    ReLU r13(.data_in(data_in[2619:2600]), .data_out(relu_out[13]));
    ReLU r14(.data_in(data_in[2599:2580]), .data_out(relu_out[14]));
    ReLU r15(.data_in(data_in[2579:2560]), .data_out(relu_out[15]));
    ReLU r16(.data_in(data_in[2559:2540]), .data_out(relu_out[16]));
    ReLU r17(.data_in(data_in[2539:2520]), .data_out(relu_out[17]));
    ReLU r18(.data_in(data_in[2519:2500]), .data_out(relu_out[18]));
    ReLU r19(.data_in(data_in[2499:2480]), .data_out(relu_out[19]));
    ReLU r20(.data_in(data_in[2479:2460]), .data_out(relu_out[20]));
    ReLU r21(.data_in(data_in[2459:2440]), .data_out(relu_out[21]));
    ReLU r22(.data_in(data_in[2439:2420]), .data_out(relu_out[22]));
    ReLU r23(.data_in(data_in[2419:2400]), .data_out(relu_out[23]));
    ReLU r24(.data_in(data_in[2399:2380]), .data_out(relu_out[24]));
    ReLU r25(.data_in(data_in[2379:2360]), .data_out(relu_out[25]));
    ReLU r26(.data_in(data_in[2359:2340]), .data_out(relu_out[26]));
    ReLU r27(.data_in(data_in[2339:2320]), .data_out(relu_out[27]));
    ReLU r28(.data_in(data_in[2319:2300]), .data_out(relu_out[28]));
    ReLU r29(.data_in(data_in[2299:2280]), .data_out(relu_out[29]));
    ReLU r30(.data_in(data_in[2279:2260]), .data_out(relu_out[30]));
    ReLU r31(.data_in(data_in[2259:2240]), .data_out(relu_out[31]));
    ReLU r32(.data_in(data_in[2239:2220]), .data_out(relu_out[32]));
    ReLU r33(.data_in(data_in[2219:2200]), .data_out(relu_out[33]));
    ReLU r34(.data_in(data_in[2199:2180]), .data_out(relu_out[34]));
    ReLU r35(.data_in(data_in[2179:2160]), .data_out(relu_out[35]));
    ReLU r36(.data_in(data_in[2159:2140]), .data_out(relu_out[36]));
    ReLU r37(.data_in(data_in[2139:2120]), .data_out(relu_out[37]));
    ReLU r38(.data_in(data_in[2119:2100]), .data_out(relu_out[38]));
    ReLU r39(.data_in(data_in[2099:2080]), .data_out(relu_out[39]));
    ReLU r40(.data_in(data_in[2079:2060]), .data_out(relu_out[40]));
    ReLU r41(.data_in(data_in[2059:2040]), .data_out(relu_out[41]));
    ReLU r42(.data_in(data_in[2039:2020]), .data_out(relu_out[42]));
    ReLU r43(.data_in(data_in[2019:2000]), .data_out(relu_out[43]));
    ReLU r44(.data_in(data_in[1999:1980]), .data_out(relu_out[44]));
    ReLU r45(.data_in(data_in[1979:1960]), .data_out(relu_out[45]));
    ReLU r46(.data_in(data_in[1959:1940]), .data_out(relu_out[46]));
    ReLU r47(.data_in(data_in[1939:1920]), .data_out(relu_out[47]));
    ReLU r48(.data_in(data_in[1919:1900]), .data_out(relu_out[48]));
    ReLU r49(.data_in(data_in[1899:1880]), .data_out(relu_out[49]));
    ReLU r50(.data_in(data_in[1879:1860]), .data_out(relu_out[50]));
    ReLU r51(.data_in(data_in[1859:1840]), .data_out(relu_out[51]));
    ReLU r52(.data_in(data_in[1839:1820]), .data_out(relu_out[52]));
    ReLU r53(.data_in(data_in[1819:1800]), .data_out(relu_out[53]));
    ReLU r54(.data_in(data_in[1799:1780]), .data_out(relu_out[54]));
    ReLU r55(.data_in(data_in[1779:1760]), .data_out(relu_out[55]));
    ReLU r56(.data_in(data_in[1759:1740]), .data_out(relu_out[56]));
    ReLU r57(.data_in(data_in[1739:1720]), .data_out(relu_out[57]));
    ReLU r58(.data_in(data_in[1719:1700]), .data_out(relu_out[58]));
    ReLU r59(.data_in(data_in[1699:1680]), .data_out(relu_out[59]));
    ReLU r60(.data_in(data_in[1679:1660]), .data_out(relu_out[60]));
    ReLU r61(.data_in(data_in[1659:1640]), .data_out(relu_out[61]));
    ReLU r62(.data_in(data_in[1639:1620]), .data_out(relu_out[62]));
    ReLU r63(.data_in(data_in[1619:1600]), .data_out(relu_out[63]));
    ReLU r64(.data_in(data_in[1599:1580]), .data_out(relu_out[64]));
    ReLU r65(.data_in(data_in[1579:1560]), .data_out(relu_out[65]));
    ReLU r66(.data_in(data_in[1559:1540]), .data_out(relu_out[66]));
    ReLU r67(.data_in(data_in[1539:1520]), .data_out(relu_out[67]));
    ReLU r68(.data_in(data_in[1519:1500]), .data_out(relu_out[68]));
    ReLU r69(.data_in(data_in[1499:1480]), .data_out(relu_out[69]));
    ReLU r70(.data_in(data_in[1479:1460]), .data_out(relu_out[70]));
    ReLU r71(.data_in(data_in[1459:1440]), .data_out(relu_out[71]));
    ReLU r72(.data_in(data_in[1439:1420]), .data_out(relu_out[72]));
    ReLU r73(.data_in(data_in[1419:1400]), .data_out(relu_out[73]));
    ReLU r74(.data_in(data_in[1399:1380]), .data_out(relu_out[74]));
    ReLU r75(.data_in(data_in[1379:1360]), .data_out(relu_out[75]));
    ReLU r76(.data_in(data_in[1359:1340]), .data_out(relu_out[76]));
    ReLU r77(.data_in(data_in[1339:1320]), .data_out(relu_out[77]));
    ReLU r78(.data_in(data_in[1319:1300]), .data_out(relu_out[78]));
    ReLU r79(.data_in(data_in[1299:1280]), .data_out(relu_out[79]));
    ReLU r80(.data_in(data_in[1279:1260]), .data_out(relu_out[80]));
    ReLU r81(.data_in(data_in[1259:1240]), .data_out(relu_out[81]));
    ReLU r82(.data_in(data_in[1239:1220]), .data_out(relu_out[82]));
    ReLU r83(.data_in(data_in[1219:1200]), .data_out(relu_out[83]));
    ReLU r84(.data_in(data_in[1199:1180]), .data_out(relu_out[84]));
    ReLU r85(.data_in(data_in[1179:1160]), .data_out(relu_out[85]));
    ReLU r86(.data_in(data_in[1159:1140]), .data_out(relu_out[86]));
    ReLU r87(.data_in(data_in[1139:1120]), .data_out(relu_out[87]));
    ReLU r88(.data_in(data_in[1119:1100]), .data_out(relu_out[88]));
    ReLU r89(.data_in(data_in[1099:1080]), .data_out(relu_out[89]));
    ReLU r90(.data_in(data_in[1079:1060]), .data_out(relu_out[90]));
    ReLU r91(.data_in(data_in[1059:1040]), .data_out(relu_out[91]));
    ReLU r92(.data_in(data_in[1039:1020]), .data_out(relu_out[92]));
    ReLU r93(.data_in(data_in[1019:1000]), .data_out(relu_out[93]));
    ReLU r94(.data_in(data_in[999:980]), .data_out(relu_out[94]));
    ReLU r95(.data_in(data_in[979:960]), .data_out(relu_out[95]));
    ReLU r96(.data_in(data_in[959:940]), .data_out(relu_out[96]));
    ReLU r97(.data_in(data_in[939:920]), .data_out(relu_out[97]));
    ReLU r98(.data_in(data_in[919:900]), .data_out(relu_out[98]));
    ReLU r99(.data_in(data_in[899:880]), .data_out(relu_out[99]));
    ReLU r100(.data_in(data_in[879:860]), .data_out(relu_out[100]));
    ReLU r101(.data_in(data_in[859:840]), .data_out(relu_out[101]));
    ReLU r102(.data_in(data_in[839:820]), .data_out(relu_out[102]));
    ReLU r103(.data_in(data_in[819:800]), .data_out(relu_out[103]));
    ReLU r104(.data_in(data_in[799:780]), .data_out(relu_out[104]));
    ReLU r105(.data_in(data_in[779:760]), .data_out(relu_out[105]));
    ReLU r106(.data_in(data_in[759:740]), .data_out(relu_out[106]));
    ReLU r107(.data_in(data_in[739:720]), .data_out(relu_out[107]));
    ReLU r108(.data_in(data_in[719:700]), .data_out(relu_out[108]));
    ReLU r109(.data_in(data_in[699:680]), .data_out(relu_out[109]));
    ReLU r110(.data_in(data_in[679:660]), .data_out(relu_out[110]));
    ReLU r111(.data_in(data_in[659:640]), .data_out(relu_out[111]));
    ReLU r112(.data_in(data_in[639:620]), .data_out(relu_out[112]));
    ReLU r113(.data_in(data_in[619:600]), .data_out(relu_out[113]));
    ReLU r114(.data_in(data_in[599:580]), .data_out(relu_out[114]));
    ReLU r115(.data_in(data_in[579:560]), .data_out(relu_out[115]));
    ReLU r116(.data_in(data_in[559:540]), .data_out(relu_out[116]));
    ReLU r117(.data_in(data_in[539:520]), .data_out(relu_out[117]));
    ReLU r118(.data_in(data_in[519:500]), .data_out(relu_out[118]));
    ReLU r119(.data_in(data_in[499:480]), .data_out(relu_out[119]));
    ReLU r120(.data_in(data_in[479:460]), .data_out(relu_out[120]));
    ReLU r121(.data_in(data_in[459:440]), .data_out(relu_out[121]));
    ReLU r122(.data_in(data_in[439:420]), .data_out(relu_out[122]));
    ReLU r123(.data_in(data_in[419:400]), .data_out(relu_out[123]));
    ReLU r124(.data_in(data_in[399:380]), .data_out(relu_out[124]));
    ReLU r125(.data_in(data_in[379:360]), .data_out(relu_out[125]));
    ReLU r126(.data_in(data_in[359:340]), .data_out(relu_out[126]));
    ReLU r127(.data_in(data_in[339:320]), .data_out(relu_out[127]));
    ReLU r128(.data_in(data_in[319:300]), .data_out(relu_out[128]));
    ReLU r129(.data_in(data_in[299:280]), .data_out(relu_out[129]));
    ReLU r130(.data_in(data_in[279:260]), .data_out(relu_out[130]));
    ReLU r131(.data_in(data_in[259:240]), .data_out(relu_out[131]));
    ReLU r132(.data_in(data_in[239:220]), .data_out(relu_out[132]));
    ReLU r133(.data_in(data_in[219:200]), .data_out(relu_out[133]));
    ReLU r134(.data_in(data_in[199:180]), .data_out(relu_out[134]));
    ReLU r135(.data_in(data_in[179:160]), .data_out(relu_out[135]));
    ReLU r136(.data_in(data_in[159:140]), .data_out(relu_out[136]));
    ReLU r137(.data_in(data_in[139:120]), .data_out(relu_out[137]));
    ReLU r138(.data_in(data_in[119:100]), .data_out(relu_out[138]));
    ReLU r139(.data_in(data_in[99:80]), .data_out(relu_out[139]));
    ReLU r140(.data_in(data_in[79:60]), .data_out(relu_out[140]));
    ReLU r141(.data_in(data_in[59:40]), .data_out(relu_out[141]));
    ReLU r142(.data_in(data_in[39:20]), .data_out(relu_out[142]));
    ReLU r143(.data_in(data_in[19:0]), .data_out(relu_out[143]));
    
    Pooling p0(.in0(relu_out[0]), .in1(relu_out[1]), .in2(relu_out[12]), .in3(relu_out[13]), .out(pooling_out[287:280]));
    Pooling p1(.in0(relu_out[2]), .in1(relu_out[3]), .in2(relu_out[14]), .in3(relu_out[15]), .out(pooling_out[279:272]));
    Pooling p2(.in0(relu_out[4]), .in1(relu_out[5]), .in2(relu_out[16]), .in3(relu_out[17]), .out(pooling_out[271:264]));
    Pooling p3(.in0(relu_out[6]), .in1(relu_out[7]), .in2(relu_out[18]), .in3(relu_out[19]), .out(pooling_out[263:256]));
    Pooling p4(.in0(relu_out[8]), .in1(relu_out[9]), .in2(relu_out[20]), .in3(relu_out[21]), .out(pooling_out[255:248]));
    Pooling p5(.in0(relu_out[10]), .in1(relu_out[11]), .in2(relu_out[22]), .in3(relu_out[23]), .out(pooling_out[247:240]));
    Pooling p6(.in0(relu_out[24]), .in1(relu_out[25]), .in2(relu_out[36]), .in3(relu_out[37]), .out(pooling_out[239:232]));
    Pooling p7(.in0(relu_out[26]), .in1(relu_out[27]), .in2(relu_out[38]), .in3(relu_out[39]), .out(pooling_out[231:224]));
    Pooling p8(.in0(relu_out[28]), .in1(relu_out[29]), .in2(relu_out[40]), .in3(relu_out[41]), .out(pooling_out[223:216]));
    Pooling p9(.in0(relu_out[30]), .in1(relu_out[31]), .in2(relu_out[42]), .in3(relu_out[43]), .out(pooling_out[215:208]));
    Pooling p10(.in0(relu_out[32]), .in1(relu_out[33]), .in2(relu_out[44]), .in3(relu_out[45]), .out(pooling_out[207:200]));
    Pooling p11(.in0(relu_out[34]), .in1(relu_out[35]), .in2(relu_out[46]), .in3(relu_out[47]), .out(pooling_out[199:192]));
    Pooling p12(.in0(relu_out[48]), .in1(relu_out[49]), .in2(relu_out[60]), .in3(relu_out[61]), .out(pooling_out[191:184]));
    Pooling p13(.in0(relu_out[50]), .in1(relu_out[51]), .in2(relu_out[62]), .in3(relu_out[63]), .out(pooling_out[183:176]));
    Pooling p14(.in0(relu_out[52]), .in1(relu_out[53]), .in2(relu_out[64]), .in3(relu_out[65]), .out(pooling_out[175:168]));
    Pooling p15(.in0(relu_out[54]), .in1(relu_out[55]), .in2(relu_out[66]), .in3(relu_out[67]), .out(pooling_out[167:160]));
    Pooling p16(.in0(relu_out[56]), .in1(relu_out[57]), .in2(relu_out[68]), .in3(relu_out[69]), .out(pooling_out[159:152]));
    Pooling p17(.in0(relu_out[58]), .in1(relu_out[59]), .in2(relu_out[70]), .in3(relu_out[71]), .out(pooling_out[151:144]));
    Pooling p18(.in0(relu_out[72]), .in1(relu_out[73]), .in2(relu_out[84]), .in3(relu_out[85]), .out(pooling_out[143:136]));
    Pooling p19(.in0(relu_out[74]), .in1(relu_out[75]), .in2(relu_out[86]), .in3(relu_out[87]), .out(pooling_out[135:128]));
    Pooling p20(.in0(relu_out[76]), .in1(relu_out[77]), .in2(relu_out[88]), .in3(relu_out[89]), .out(pooling_out[127:120]));
    Pooling p21(.in0(relu_out[78]), .in1(relu_out[79]), .in2(relu_out[90]), .in3(relu_out[91]), .out(pooling_out[119:112]));
    Pooling p22(.in0(relu_out[80]), .in1(relu_out[81]), .in2(relu_out[92]), .in3(relu_out[93]), .out(pooling_out[111:104]));
    Pooling p23(.in0(relu_out[82]), .in1(relu_out[83]), .in2(relu_out[94]), .in3(relu_out[95]), .out(pooling_out[103:96]));
    Pooling p24(.in0(relu_out[96]), .in1(relu_out[97]), .in2(relu_out[108]), .in3(relu_out[109]), .out(pooling_out[95:88]));
    Pooling p25(.in0(relu_out[98]), .in1(relu_out[99]), .in2(relu_out[110]), .in3(relu_out[111]), .out(pooling_out[87:80]));
    Pooling p26(.in0(relu_out[100]), .in1(relu_out[101]), .in2(relu_out[112]), .in3(relu_out[113]), .out(pooling_out[79:72]));
    Pooling p27(.in0(relu_out[102]), .in1(relu_out[103]), .in2(relu_out[114]), .in3(relu_out[115]), .out(pooling_out[71:64]));
    Pooling p28(.in0(relu_out[104]), .in1(relu_out[105]), .in2(relu_out[116]), .in3(relu_out[117]), .out(pooling_out[63:56]));
    Pooling p29(.in0(relu_out[106]), .in1(relu_out[107]), .in2(relu_out[118]), .in3(relu_out[119]), .out(pooling_out[55:48]));
    Pooling p30(.in0(relu_out[120]), .in1(relu_out[121]), .in2(relu_out[132]), .in3(relu_out[133]), .out(pooling_out[47:40]));
    Pooling p31(.in0(relu_out[122]), .in1(relu_out[123]), .in2(relu_out[134]), .in3(relu_out[135]), .out(pooling_out[39:32]));
    Pooling p32(.in0(relu_out[124]), .in1(relu_out[125]), .in2(relu_out[136]), .in3(relu_out[137]), .out(pooling_out[31:24]));
    Pooling p33(.in0(relu_out[126]), .in1(relu_out[127]), .in2(relu_out[138]), .in3(relu_out[139]), .out(pooling_out[23:16]));
    Pooling p34(.in0(relu_out[128]), .in1(relu_out[129]), .in2(relu_out[140]), .in3(relu_out[141]), .out(pooling_out[15:8]));
    Pooling p35(.in0(relu_out[130]), .in1(relu_out[131]), .in2(relu_out[142]), .in3(relu_out[143]), .out(pooling_out[7:0]));
        
    CSR_encoder csr1(.data_in(pooling_out), .enable(en_encoder), .clk(clk), .row_size(row_size), .index_pointer(index_pointer), .row(row), .data(data), .store(store), .done(done));
    
    assign out_port = (en_pooling == 1)? 0: {relu_out[0],relu_out[1],relu_out[12],relu_out[13]};

endmodule