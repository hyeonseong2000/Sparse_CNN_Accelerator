// ROMs Using Block RAM Resources.
// File: rams_sp_rom_1.v
//
module weight_index_ROM (clk, en, addr, rout);
    input clk;
    input en;
    input [6:0] addr;
    output [47:0] rout;

(*rom_style = "block" *) reg [47:0] rowptr;

    always @(posedge clk) begin
        if (en)
            case(addr)
            7'd0: rowptr <= 48'b000000000000000100000100000001000000010100000110;
            7'd1: rowptr <= 48'b000000000000000000000000000000100000001100000011;
            7'd2: rowptr <= 48'b000000000000000100000001000000010000000100000001;
            7'd3: rowptr <= 48'b000000000000000100000010000000100000011100001000;
            7'd4: rowptr <= 48'b000000000000000100000010000000110000011000000110;
            7'd5: rowptr <= 48'b000000000000000000000000000000100000010000001000;
            7'd6: rowptr <= 48'b000000000000000000000000000000000000000000000001;
            7'd7: rowptr <= 48'b000000000000000000000000000000010000001000000010;
            7'd8: rowptr <= 48'b000000000000001000000100000001110000100000001000;
            7'd9: rowptr <= 48'b000000000000000000000001000000010000001100000100;
            7'd10: rowptr <= 48'b000000000000000000000010000000110000010000000100;
            7'd11: rowptr <= 48'b000000000000000100000010000000110000001100000100;
            7'd12: rowptr <= 48'b000000000000000100000011000001000000010100000110;
            7'd13: rowptr <= 48'b000000000000001000000011000001000000010100000101;
            7'd14: rowptr <= 48'b000000000000000100000011000001010000100000001001;
            7'd15: rowptr <= 48'b000000000000010000000110000001110000011100001000;
            7'd16: rowptr <= 48'b000000000000000100000011000001100000011100001000;
            7'd17: rowptr <= 48'b000000000000001100000110000001110000011100001000;
            7'd18: rowptr <= 48'b000000000000000100000001000000100000001000000011;
            7'd19: rowptr <= 48'b000000000000000100000011000000110000010000000110;
            7'd20: rowptr <= 48'b000000000000000100000010000001000000010100000101;
            7'd21: rowptr <= 48'b000000000000000000000000000000010000000100000011;
            7'd22: rowptr <= 48'b000000000000001000000100000001100000100000001000;
            7'd23: rowptr <= 48'b000000000000000000000000000000000000000000000011;
            7'd24: rowptr <= 48'b000000000000001000000010000000100000001000000010;
            7'd25: rowptr <= 48'b000000000000001100000101000001100000100000001010;
            7'd26: rowptr <= 48'b000000000000001000000100000001100000100000001001;
            7'd27: rowptr <= 48'b000000000000000100000011000000110000001100000100;
            7'd28: rowptr <= 48'b000000000000001100000110000010000000100100001011;
            7'd29: rowptr <= 48'b000000000000001100000011000000110000001100000011;
            7'd30: rowptr <= 48'b000000000000000100000001000000010000000100000010;
            7'd31: rowptr <= 48'b000000000000000100000010000000100000001000000010;
            7'd32: rowptr <= 48'b000000000000000000000001000000100000001000000011;
            7'd33: rowptr <= 48'b000000000000000100000011000001000000010100000101;
            7'd34: rowptr <= 48'b000000000000001000000110000001110000100100001010;
            7'd35: rowptr <= 48'b000000000000000000000001000000100000001000000100;
            7'd36: rowptr <= 48'b000000000000000000000000000000100000001100000101;
            7'd37: rowptr <= 48'b000000000000001000000010000000110000010000000110;
            7'd38: rowptr <= 48'b000000000000000100000011000001010000010100000101;
            7'd39: rowptr <= 48'b000000000000001000000010000001000000010100001000;
            7'd40: rowptr <= 48'b000000000000000000000001000000110000010000000110;
            7'd41: rowptr <= 48'b000000000000000100000010000000110000001100000101;
            7'd42: rowptr <= 48'b000000000000001000000100000001000000010000000100;
            7'd43: rowptr <= 48'b000000000000010100000101000001010000010100000111;
            7'd44: rowptr <= 48'b000000000000000000000010000001000000011000000110;
            7'd45: rowptr <= 48'b000000000000001100000100000001010000011100001001;
            7'd46: rowptr <= 48'b000000000000000000000000000000010000000100000010;
            7'd47: rowptr <= 48'b000000000000000000000000000000100000010000000110;
            7'd48: rowptr <= 48'b000000000000001000000011000001000000010000000100;
            7'd49: rowptr <= 48'b000000000000000000000001000000010000001000000100;
            7'd50: rowptr <= 48'b000000000000000000000010000001000000011100001001;
            7'd51: rowptr <= 48'b000000000000001000000100000001010000010100000110;
            7'd52: rowptr <= 48'b000000000000000000000000000000100000001100000100;
            7'd53: rowptr <= 48'b000000000000001000000010000000100000010100000101;
            7'd54: rowptr <= 48'b000000000000000100000001000000100000001100000100;
            7'd55: rowptr <= 48'b000000000000000100000010000001000000010000000110;
            7'd56: rowptr <= 48'b000000000000001000000100000001100000011100001000;
            7'd57: rowptr <= 48'b000000000000000000000000000000000000001000000011;
            7'd58: rowptr <= 48'b000000000000000000000011000001110000101000001011;
            7'd59: rowptr <= 48'b000000000000000100000100000001010000011100001000;
            7'd60: rowptr <= 48'b000000000000001000000010000000100000001100000011;
            7'd61: rowptr <= 48'b000000000000000100000100000001000000010000000101;
            7'd62: rowptr <= 48'b000000000000001000000011000001000000100000001001;
            7'd63: rowptr <= 48'b000000000000001000000011000001000000010100000111;
            7'd64: rowptr <= 48'b000000000000000000000010000000110000010100000101;
            7'd65: rowptr <= 48'b000000000000000000000010000001000000010000000111;
            7'd66: rowptr <= 48'b000000000000001000000010000001000000010100000110;
            7'd67: rowptr <= 48'b000000000000000100000001000000100000001100000100;
            7'd68: rowptr <= 48'b000000000000001100000100000001010000011000001000;
            7'd69: rowptr <= 48'b000000000000000100000010000000100000001100000100;
            7'd70: rowptr <= 48'b000000000000000100000001000000010000001100000011;
            7'd71: rowptr <= 48'b000000000000001000000010000000110000001100000100;
            7'd72: rowptr <= 48'b000000000000000100000010000000110000010100000110;
            7'd73: rowptr <= 48'b000000000000000100000010000001000000011000000110;
            7'd74: rowptr <= 48'b000000000000000000000000000000100000001100000100;
            7'd75: rowptr <= 48'b000000000000000100000011000001000000010100000110;
            7'd76: rowptr <= 48'b000000000000000000000011000000110000001100000011;
            7'd77: rowptr <= 48'b000000000000000000000001000000100000001100000011;
            7'd78: rowptr <= 48'b000000000000001000000011000001010000010100000110;
            7'd79: rowptr <= 48'b000000000000001000000011000001010000011000000110;
            7'd80: rowptr <= 48'b000000000000000000000001000000110000010000000101;
            7'd81: rowptr <= 48'b000000000000000100000010000000110000010000000100;
            7'd82: rowptr <= 48'b000000000000000100000001000001000000010000000100;
            7'd83: rowptr <= 48'b000000000000000100000010000000100000001100000011;
            7'd84: rowptr <= 48'b000000000000000000000000000000000000000100000001;
            7'd85: rowptr <= 48'b000000000000000000000000000000000000001000000100;
            7'd86: rowptr <= 48'b000000000000000000000001000000010000001100000100;
            7'd87: rowptr <= 48'b000000000000000100000001000000100000010000000100;
            7'd88: rowptr <= 48'b000000000000001000000011000001010000010100000111;
            7'd89: rowptr <= 48'b000000000000000100000001000000010000001000000011;
            7'd90: rowptr <= 48'b00000000_00000001_00000001_00000001_00000001_00000001;
            7'd91: rowptr <= 48'b000000000000000100000010000000110000010000000101;
            7'd92: rowptr <= 48'b000000000000001100000101000001110000100000001010;
            7'd93: rowptr <= 48'b000000000000000000000010000000110000010000000100;
            7'd94: rowptr <= 48'b000000000000000000000000000000100000001100000111;
            7'd95: rowptr <= 48'b000000000000001100000100000001000000010100000101;
            7'd96: rowptr <= 48'b000000000000000100000010000000100000010000000101;
            7'd97: rowptr <= 48'b000000000000000000000000000000000000000100000010;
            7'd98: rowptr <= 48'b000000000000000000000001000000100000001000000011;
            7'd99: rowptr <= 48'b000000000000001100000011000001000000010100000110;
            7'd100: rowptr <= 48'b000000000000000000000000000000010000001000000011;
            7'd101: rowptr <= 48'b000000000000000000000010000000110000010000000101;
            endcase
    end

    assign rout = rowptr;

endmodule